module alu(
	input [31:0] dataA, dataBi,
	
)
